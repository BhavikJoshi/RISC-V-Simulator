module reorder_buffer ();

endmodule